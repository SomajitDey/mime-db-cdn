application/x-virtualbox-vhd
